Colpitt oscillator using BJT

.MODEL QBC547BP NPN(IS=1.8E-14 BF=400 NF=0.9955 VAF=80 IKF=0.14 
+ ISE=5E-14 NE=1.46 BR=35.5 NR=1.005 VAR=12.5 IKR=0.03 ISC=1.72E-13 
+ NC=1.27 RB=0.56 RE=0.6 RC=0.25 CJE=1.3E-11 TF=6.4E-10 CJC=4E-12 VJC=0.54 TR=5.072E-8 )

Vcc 2 0 dc 9V
R1 2 1 100k
R2 1 0 5k
R3 2 3 1k
R4 6 0 10k

Q1 3 1 6 QBC547BP

C3 5 1 100pf
c1 5 0 0.01uf
C2 0 4 0.01uf
C4 6 0 100nf
C5 3 4 100pf

L1 5 4 10mh

.control
tran 0.1us 500u 200u UIC
run
set color0 = white
set control = black
plot V(4)
.endc
.end
Active bandpass filter

.include LF356.MOD
XU1 3 2 7 4 6 LF356/NS
XU2 13 12 17 14 16 LF356/NS

Vin 1 0 AC 1 DC 0 
V7 7 0 12V
V4 4 0 -12V
V17 17 0 12V
V14 14 0 -12V
R1 3 0 1K
R2 2 0 100k
R3 2 6 1K
R4 6 13 10K
R5 12 0 1K
R6 12 16 1K
R7 16 0 1
C1 1 3 10uF 
C2 13 0 1pF

.ac dec 10 1 80Meg
.control
run
set color0 = white
set color1 = black
set color2 = blue
set Xbrushwidth = 2
plot v(16)

.endc
.end
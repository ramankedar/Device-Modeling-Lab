Integrator using op-amp

.INCLUDE LF356.MOD
XU1 1 0 6 5 3 LF356/NS

Vin 2 0 SIN(0 10 50)
R1 2 1 10k
C1 1 3 100nF
R2 1 3 2.2M
V2 0 6 dc 10
V3 5 0 dc 10

.control
tran 1us 0.1s
*set Xbrushwidth = 2
run
set color0 = white
set color1 = black
plot V(2) V(3)

.endc
.end

NOT Gate

vdd 3 0 dc 5v

m1 3 1 2 3 mos1 l=10u w=100u
.model mos1 pmos vto=1.5v kp=200u

m2 2 1 0 0 mos2 l=10u w=100u
.model mos2 nmos vto=1.5v kp=200u

vin 1 0 pulse(0 5 0 0 100ns 800ns)

.tran 10ns 1200ns
.control
run
plot v(1) v(2)

.endc
.end
N-channel Mosfet characteristics

v1 2 0 5
v2 1 0 1
r1 2 3 0
r2 1 4 0
m1 3 4 0 0 NFET

.model NFET NMOS

.dc v1 0 3 1m
.options savecurrents
.control
run

set color0 = white
set color1 = black
set color2 = red

plot @r1[i]

.endc
.end
XOR USING NAND

V1 1 0 PULSE(0 5 0 0 0 10ms 20ms)
V2 2 0 PULSE(0 5 0 0 0 20ms 40ms)
X1 1 2 3 NAND
X2 1 3 4 NAND
X3 2 3 5 NAND
X4 4 5 Y NAND

.SUBCKT NAND 1 2 Y
D1 M 1 D
D2 M 2 D
D3 M 21 D
Q1 Y 21 0 BJT1
R1 V M 80K
R2 V Y 80K
V1 V 0 5
.model D D
.MODEL BJT1 NPN(BF=150 CJC=10pf CJE=10pf IS=1E-16 RE=1k RC=1k RB=1k)
.ENDS
.CONTROL
TRAN 0.01ms 80ms
PLOT v(1)+30 v(2)+15 v(Y)

.ENDC
.END
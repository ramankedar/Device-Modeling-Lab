Active bandstop filter

.include LF356.MOD
XU1 3 2 7 4 6 LF356/NS
XU2 13 12 17 14 16 LF356/NS
XU3 23 22 27 24 26 LF356/NS

Vin 1 0 AC 1 DC 0 
V17 7 0 12V
V14 4 0 -12V
V27 17 0 12V
V24 14 0 -12V
V37 27 0 12V
V34 34 0 -12V

R1 1 3 10k
C1 3 0 1uF
C2 1 13 1nF
R2 13 0 10k
R3 6 32 1k
R4 16 32 1k
R5 32 36 1k

.ac dec 100 1 1Meg
.control
run
set color0 = white
set color1 = black
set color2 = blue
set Xbrushwidth = 2
plot V(36)

.endc
.end

Full Wave Rectifier with Resistance as a Load

vin 0 1 sin(0 2 75 0 0 0)
D1 2 1 D1N4148
D2 1 3 D1N4148
D3 0 3 D1N4148
D4 2 0 D1N4148
R 3 2 10k

.model D1N4148 D (IS=0.1PA, RS=16 CJO=2PF TT=12N BV=100 IBV=0.1PA)                                            
.TRAN 1u 40m
.CONTROL
run
set color0 = white
set color1 = black
PLOT V(3)-V(2) V(1)
*PLOT I(3) I(1)
PLOT (V(3)-V(2))/10k

.ENDC
.END
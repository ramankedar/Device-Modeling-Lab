NAND gate using CMOS

vdd 1 0 dc 5v

m1 1 2 4 1 mos1 l=10u w=100u
.model mos1 pmos vto=1.5v kp=200u

m2 1 3 4 1 mos2 l=10u w=100u
.model mos2 pmos vto=1.5v kp=200u

m3 4 2 5 5 mos3 l=10u w=100u
.model mos3 nmos vto=1.5v kp=200u

m4 5 3 0 0 mos4 l=10u w=100u
.model mos4 nmos vto=1.5v kp=200u

vin1 2 0 pulse(0 5 0 0 100ns 800ns)
vin2 3 0 pulse(5 0 0 0 100ns 800ns)

.tran 10ns 1200ns
.control
run
plot v(4) v(2) v(3)

.endc
.end
Full Wave Rectifier

V1 n0 0 SIN(0 20 1kHz)
D1 n1 n0 D
D2 n1 0 D
D3 0 n3 D
D4 n0 n3 D
R1 n3 n1 1k

.model D D

.CONTROL 
TRAN 0.02ms 20ms 
PLOT V(n1) V(0)

.ENDC a
.END
Common Drain Amplifier using JFET

vin 1 0 sine(0 5m 100 0 0 0)
c1 1 2 10u
v2 3 0 15
r2 4 0 10k
c2 4 5 10u
rL 5 0 10K

J1 3 2 4 NJF

.model NJF NJF
.tran 1u 20m
.control
run
set color0=white
set color1=black
set color2=green
set color3=red
set color4=blue
set Xbrushwidth=2
plot v(1) v(5)

.endc
.end
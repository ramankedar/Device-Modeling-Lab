A simple RC High Pass Filter 

V1 n0 0 SIN(0 10 1kHz)
C1 n0 n1 3.3nF
R1 n1 0 1k

.CONTROL 
TRAN 0.01ms 10ms 
PLOT V(n0) V(n1)

.ENDC 
.END
Non-inverting summer

.INCLUDE UA741.MOD
XU1 0 2 7 4 6 UA741

V1 1 0 SIN(0 5 1kHz)
V2 2 0 SIN(0 5 1kHz)
V7 7 0 12V
V4 4 0 -12V
R1 1 3 1K
R2 2 3 1K
R3 3 6 10K

.tran 1us 0.01s
.control
run

set color0 = white
set color1 = black
set Xbrushwidth = 2
plot V(1)+10 V(3)+5 V(6)/2-7
.endc
.end

3 INPUT AND GATE USING NAND

VA 1 0 PULSE(0 5 0 0 0 10ms 20ms)
VB 2 0 PULSE(0 5 0 0 0 20ms 40ms)
VC 3 0 PULSE(0 5 0 0 0 30ms 60ms)
X1 1 2 4 NAND
X2 4 4 6 NAND
X3 6 3 Z NAND
X4 Z Z Y NAND
* SUBCKT NAND GATE
.SUBCKT NAND 1 2 Y
D2 M 2 D
D1 M 1 D
D3 M 21 D
Q1 Y 21 0 BJT1
R1 V M 80K
R2 V Y 80K
V1 V 0 5
.model D D
.MODEL BJT1 NPN(BF=150 CJC=10pf CJE=10pf IS=1E-16 RE=1k RC=1k RB=1k)
.ENDS
.CONTROL
TRAN 0.01ms 100ms
PLOT v(1)+45 v(2)+30 v(3)+15 v(Y)
.ENDC
.END

Hartley oscillator using BJT

.MODEL QBC547BP NPN(IS=1.8E-14 BF=400 NF=0.9955 VAF=80 IKF=0.14 
+ ISE=5E-14 NE=1.46 BR=35.5 NR=1.005 VAR=12.5 IKR=0.03 ISC=1.72E-13 
+ NC=1.27 RB=0.56 RE=0.6 RC=0.25 CJE=1.3E-11 TF=6.4E-10 CJC=4E-12 
+ VJC=0.54 TR=5.072E-8 )

Vcc vin 0 dc 9
R1 vin a 100k
R2 a 0 5k
R3 vin b 1k
R4 c 0 10k

Q1 a b c QBC547BP

C1 a d 100pf
C2 d out 10pf
C3 c 0 100pf
C4 b out 100pf

L1 d 0 10mh
L2 0 out 20mh

.control
tran 0.1u 500u
run
set color0 = white
set control = black
plot V(out)
.endc
.end
Positive Clipper: Negative Bias

V1 0 n1 sin(0 1 50)
D1 n2 n1 D
R1 n2 n3 100k
vol n3 0 -0.3

.model D D

.CONTROL
TRAN 0.01ms 70ms
set color0 = white
set color1 = black
PLOT V(n1) V(n2)

.ENDC
.END
Full Wave Rectifier


V1 n0 n2 SIN(0 10 1kHz)
D1 0 n0 D
D2 0 n2 D
D3 n0 n1 D
D4 n2 n1 D
R1 n1 0 1k

.model D D

.CONTROL 
TRAN 0.01ms 10ms 
PLOT V(n0)  V(n1)



.ENDC 
.END
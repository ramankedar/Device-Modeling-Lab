Edge triggering D-flip flop

.SUBCKT NAND in1 in2 out VDD
M1 out in2 Vdd Vdd p1 W=7.5u L=0.35u pd=13.5u ad=22.5p ps=13.5u as=22.5p
M2 net.1 in2 0 0 n1   W=3u   L=0.35u pd=9u    ad=9p    ps=9u    as=9p
M3 out in1 Vdd Vdd p1 W=7.5u L=0.35u pd=13.5u ad=22.5p ps=13.5u as=22.5p
M4 out in1 net.1 0 n1 W=3u   L=0.35u pd=9u    ad=9p    ps=9u    as=9p
.ENDS NAND

vcc 1 0 dc 5
v1 in1 0 pulse(0 5 0 0 0 15ms 30ms)
v2 cl 0 pulse(0 5 0 0 0 5ms 10ms)
.model n1 nmos level=49 version=3.3.0
.model p1 pmos level=49 version=3.3.0

X1 cl cl 2 1 NAND
X2 in1 2 3 1 NAND
X3 2 3 4 1 NAND
X4 2 2 5 1 NAND
X5 3 6 7 1 NAND
X6 4 7 6 1 NAND
X7 7 5 8 1 NAND
X8 8 5 9 1 NAND
X9 9 op 10 1 NAND
X10 8 10 op 1 NAND

.control
tran 0.01m 100m
set color0=white
set color1=black
set color2=blue
set color3=green
set color4=red
set xbrushwidth=2
plot v(op),v(cl)+6,v(in1)+15

.endc
.end
Clamper circuit

V1 n0 0 sin(0 25 1KHz)
C1 n0 n1 10uF
R1 n1 o 1k
D1 0 n1 D

.model D D

.CONTROL
TRAN 0.01ms 5ms
set color0 = white
set color1 = black
PLOT V(n0) V(n1)

.ENDC
.END